module RV32IA(inst,PC_out,clk_in,enable,inst_fetc,reset);

input [31:0] inst;//inst(instruction to drive the cpu)
input clk_in,enable,reset;
output[31:0] PC_out;
output inst_fetc;
logic [31:0] PC;
logic [3:0] operation;//operation({func_7 merge with forced signed "1", funct_3[2:0]})
logic [1:0] ALUop,WB_Mux_sel,ALU_SRC_B;//ALUop( to use as the indicator for the ALU_control to decide what would happen to the ALU outside the ALU instructions)
logic [6:0] opcode;//opcode(operation code field)
logic [31:0]ALU_out,ALU_out_Latched,ALU_in_rs1_Latched,ALU_in_rs2_Latched,
				imm,
				imm_out,imm_out_latched,
				MUX_OUT,
				Write_Data_mem,
				Read_Data_mem,
				complete_Read_Data_mem;//ALU_out(the result calculated by the integer ALU),imm(the immediate value generated by imm_gen module)

logic [31:0]ALU_in_rs1,
				ALU_in_rs2,
				ALU_SRC_B_MUX,
				ALU_SRC_A_MUX;//ALU_in_rs1(read the value from register 1 then wired to the A port of the ALU),ALU_in_rs2(read the value from register 2 then wired to the B port of the ALU)

logic [4:0] RS1,
				RS2,
				RSD;

logic clr,
		Reg_Write,
		Mem_Write,
		Mem_Read,
		ALU_SRC_A,
		PC_Write,
		more,even,less,
		done,
		Debug,Debug_signal,clk;

///* test 

	ALU_control ALU_ctrl(
								.opcode(inst[6:0]),
								.funct_7(inst[31:25]),
								.funct_3(inst[14:12]),
								.ALUop(ALUop),
								.operation(operation)
								);		
	

	
	ALU ALU(
				.result(ALU_out),
				.operation(operation),
				.a(ALU_SRC_A_MUX),
				.b(ALU_SRC_B_MUX),
				.More(more),
				.Even(even),
				.Less(less)
				);				

	Reg_32bit ALU_OUT_register(
									.enable(1'b1),
									.choose(1'b1),
									.clr(clr),
									.clk(clk),
									.Data_in(ALU_out),
									.Data_out(ALU_out_Latched)// (current PC) 
									);	
	MUX4 ALU_src_B_MUX(
						.sel(ALU_SRC_B),
						.in1(ALU_in_rs2_Latched),
						.in2(32'h4),
						.in3(imm),
						.in4(imm_out_latched),
						.MUX_OUT(ALU_SRC_B_MUX)
						);
	MUX2 ALU_src_A_MUX(
							.sel(ALU_SRC_A),
							.in1(PC),
							.in2(ALU_in_rs1_Latched),
							.out(ALU_SRC_A_MUX)
						);			
						
	Reg_32bit PC_register(
									.enable(1'b1),
									.choose(1'b1),
									.clr(clr|Debug_signal),
									.clk(PC_Write),
									.Data_in(ALU_out),
									.Data_out(PC)// (current PC) 
									);	
	//assign clock_ctrl = ~Debug_signal?PC_Write:1'b0;
	
	assign PC_out = PC;
									
	Initializer Init(.clk(clk),.enable(enable),.Debug(Debug_signal),.clr(clr),.reset(reset));//Initializing the cpu, or halting/return the cpu to debug mode.
									
	Register_file Reg_file(
									.RS1(RS1),
									.RS2(RS2),
									.RSD(RSD),
									.Data_in(MUX_OUT),
									.clr(clr),
									.Reg_Write(Reg_Write),
									.RD1(ALU_in_rs1),
									.RD2(ALU_in_rs2)
									);		

	Reg_32bit ALU_in_rs1_register(
									.enable(1'b1),
									.choose(1'b1),
									.clr(clr),
									.clk(clk),
									.Data_in(ALU_in_rs1),
									.Data_out(ALU_in_rs1_Latched)// (current PC) 
									);
	Reg_32bit ALU_in_rs2_register(
									.enable(1'b1),
									.choose(1'b1),
									.clr(clr),
									.clk(clk),
									.Data_in(ALU_in_rs2),
									.Data_out(ALU_in_rs2_Latched)// (current PC) 
									);			
	
	MUX4  			WBMUX(	.sel(WB_Mux_sel),// write back to register
									.in1(ALU_out_Latched),
									.in2(imm),
									.in3(complete_Read_Data_mem),
									.in4(),
									.MUX_OUT(MUX_OUT)
									);

	imm_gen IMM_GEN(
						.inst(inst[31:0]),
						.result(imm)
						);
	
	branch Br(
					.funct_3(inst[14:12]),
					.more(more),
					.even(even),
					.less(less),
					.imm_in(imm),
					.imm_out(imm_out)
				);

	Reg_32bit Branch_imm(
									.enable(1'b1),
									.choose(1'b1),
									.clr(clr),
									.clk(clk),
									.Data_in(imm_out),
									.Data_out(imm_out_latched)// (current PC) 
									);

	instruction_decoder inst_decode(
												.inst(inst),
												.opcode(opcode),
												.RS1(RS1),
												.RS2(RS2),
												.RSD(RSD)
												);			
												
	

	control ctrl(
						.opcode(inst[6:0]),
						.ebreak(inst[31:20]),
						.WB_Mux_sel(WB_Mux_sel),
						.ALUop(ALUop),
						.ALU_src_A(ALU_SRC_A),
						.ALU_src_B(ALU_SRC_B),
						.Reg_Write(Reg_Write),
						.Mem_Read(Mem_Read),
						.Mem_Write(Mem_Write),
						.PC_Write(PC_Write),
						.clk(clk),//problem not fix here(suggestion should add a latch to be able to unlatch the Debug )
						.Debug(Debug),
						.reset(clr|Debug_signal),//problem not fix here(suggestion should add a latch to be able to unlatch the Debug )
						.done(done)
						);
	
	assign clk = clk_in|Debug_signal;//block clk signal when Debug is raised
	
	//assign 
	///*
	always @(*)
	begin
		if(enable) Debug_signal <= Debug;
		else Debug_signal <= 'h0;
	end
	//*/
	assign inst_fetc = done & enable ;// done is when control unit is at state=0, enable is when the reset is on

	Data_Memory DMEM(
							.Write_Data(Write_Data_mem),
							.Address(ALU_out_Latched),
							.Mem_Read(Mem_Read),
							.Mem_Write(Mem_Write),
							.Read_Data(Read_Data_mem)
							);
	LD_ST_data_complete data_Read_Write_converter(
																	.opcode(inst[6:0]),
																	.funct_3(inst[14:12]),
																	.Read_Data_mem(Read_Data_mem),
																	.Write_Data_mem(ALU_in_rs2),
																	.complete_Read_Data_mem(complete_Read_Data_mem),
																	.complete_Write_Data_mem(Write_Data_mem)
																	);
//*/
		

endmodule 

//======================================================
//======================================================	
module MUX2(sel,in1,in2,out);
input sel;
input [31:0] in1,in2;
output[31:0] out;

generate
		genvar i;
	for(i=0;i<32;i++)begin : mux2
			assign out[i] = sel? in2[i]:in1[i];
	end
endgenerate

endmodule 
//======================================================
//======================================================
module MUX2_5bits(sel,in1,in2,out);
input sel;
input [4:0] in1,in2;
output[4:0] out;

	generate
			genvar i;
		for(i=0;i<5;i++)begin : mux2_5bits
				assign out[i] = sel? in2[i]:in1[i];
		end
	endgenerate

endmodule 
//======================================================
//======================================================
module Initializer(clk,enable,Debug,clr,reset);
	input enable,clk,Debug,reset;
	logic DO,latch_data;
	output clr;
	//we exploit the register characteristic of initial rising edge when clr is set to "0" the 'DO' get reset to "0"  
	//then clk rising edge update the DO to "0"
	///*
		Reg_1bit REG(
						.clr(1'b0),
						.clk(clk),
						.Data_in(1'b1),
						.Data_out(DO)
						);
	//*/
	always @(*)
	begin
			latch_data = enable; //enable=1 is clr,=0 is not clr, Debug=1 is clr,=0 is not clr  
	end
	assign clr = (latch_data ^ DO);

endmodule 

